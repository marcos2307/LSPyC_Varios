module decoder(
    input clk,
    input [4:0] in,
    output reg [17:0] out
    );



   always @(posedge clk)
        case (in)
             1  : out <= 18'b001100001100000011; //+1
             2  : out <= 18'b000011000011001100; //-1
             3  : out <= 18'b110000110000001100; //+2
             4  : out <= 18'b001100001100110000; //-2
             5  : out <= 18'b000011000011110000; //+3
             6  : out <= 18'b110000110000000011; //-3
             7  : out <= 18'b001100000011001100; //+4
             8  : out <= 18'b000011001100000011; //-4
             9  : out <= 18'b110000001100110000; //+5
            10  : out <= 18'b001100110000001100; //-5
            11  : out <= 18'b000011110000000011; //+6
            12  : out <= 18'b110000000011110000; //-6
            13  : out <= 18'b000011001100001100; //+7
            14  : out <= 18'b001100000011000011; //-7
            15  : out <= 18'b001100110000110000; //+8
            16  : out <= 18'b110000001100001100; //-8
            17  : out <= 18'b110000000011000011; //+9
            18  : out <= 18'b000011110000110000; //-9
            19  : out <= 18'b000011000011000011; //0a
            20  : out <= 18'b001100001100001100; //0b
            21  : out <= 18'b110000110000110000; //0c
            22  : out <= 18'b110000001100000011; //r
            23  : out <= 18'b001100000011110000;
            24  : out <= 18'b000011110000001100;
            25  : out <= 18'b001100110000000011;
            26  : out <= 18'b110000000011001100;
            27  : out <= 18'b000011001100110000;
        default : out <= 18'b000000000000000000;
         endcase
endmodule
